`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/05/2020 12:59:36 PM
// Design Name: 
// Module Name: errorDetect_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module recordMeta_tb();

    logic clk;
	logic resetN;
	logic dIn;
	logic samplePulse;
	logic enable;
    logic save;
    logic calc;
    logic [31:0] sig;
    logic true;
    logic complete;
    logic ready;
    logic pulseWrite;

	
    recordMaster dut(.clk, .resetN, .dIn, .samplePulse, .enable, .writeOut(save), .determineOW(calc), .owTrue(true), .complete, .owReady(ready),
        .pulseWrite, .playbackOut(sig));

	
	//Initial values
	
	initial begin
	   clk = 1;
	   resetN = 1;
       samplePulse = 1;
	   dIn = 0;
	   enable = 0;
       save = 0;
       calc = 0;
	end
	
	always begin
	   #2.5 clk = !clk;
	end

    always begin
        #5 samplePulse = !samplePulse;
    end
	
	task bitZero();
        begin
            dIn = 0;
            #10;
        end
    endtask
    task bitOne();
        begin
            dIn = 1;
            #10;
        end
    endtask
    
    task bigData();
        begin
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
        bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
        bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
        end
    endtask

    task calcSignalPassEasy();
        begin
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
        end
    endtask

    task calcSignalPassHard();
        begin
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
        end
    endtask

    task calcSignalPassEdge();
        begin
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
        end
    endtask


    task calcSignalFail();
        begin
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
        end
    endtask
    
    initial begin
        #25;
        resetN = 0;
        #45;
        resetN = 1;
        #25
        enable = 1;
        save = 1;
        #10;
        bigData();
        enable = 0;
        #10;
        wait(complete == 1);
        save = 0;
        #250;
        resetN = 0;
        #45;
        resetN = 1;
        #25
        enable = 1;
        calc = 1;
        #10;
        calcSignalPassEasy();
        enable = 0;
        #10;
        wait(complete == 1);
        #200;
        calc = 0;
        #250;
        resetN = 0;
        #45;
        resetN = 1;
        #25
        enable = 1;
        calc = 1;
        #10;
        calcSignalPassHard();
        enable = 0;
        #10;
        wait(complete == 1);
        #200;
        calc = 0;
        #250;
        resetN = 0;
        #45;
        resetN = 1;
        #25
        enable = 1;
        calc = 1;
        #10;
        calcSignalPassEdge();
        #10;
        enable = 0;
        #10;
        wait(complete == 1);
        #200;
        calc = 0;
        #250;
        resetN = 0;
        #45;
        resetN = 1;
        #25
        enable = 1;
        calc = 1;
        #10;
        calcSignalFail();
        enable = 0;
        #10;
        wait(complete == 1);
        #200;
        calc = 0;
        #250;
        $stop;
        
    end
    

endmodule
