//Part 1

in = 1;
#2000;
in = 0;
#200