`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/05/2020 12:59:36 PM
// Design Name: 
// Module Name: errorDetect_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module sigRecord_tb();

    logic clk;
	logic resetN;
	logic dIn;
	logic samplePulse; //Since we are in the early bit, this gets pulsed three times. Make sure to read the value after the third pulse
	logic enable;
    logic [31:0] sig;
    logic valid;
    logic [31:0] runningTotal;
    logic [5:0] incrementer;
    logic [8:0] baseAddr;
    logic [8:0] numFetches;
    logic enableStore;
    logic returnToBaseAddr;
    logic request;
    logic incrementAddr;
    logic [31:0] currOut;
    logic writeDBG;
    logic [7:0] pointerDBG;
	
	recordUnit rU(.clk, .resetN, .dIn, .samplePulse, .enable, .recordedOut(sig), .dataValid(valid), .runningTotal, .incrementer);
    sigStorage dut(.clk, .resetN, .baseAddr, .numFetches, .storeConfig(enableStore), .bramIn(sig), .fetch(valid), .returnToBaseAddr, .request(request), .incrementAddr, .playbackOut(currOut), .writeDBG, .pointerDBG);
    
	
	//Initial values
	
	initial begin
	   clk = 1;
	   resetN = 1;
       samplePulse = 1;
	   dIn = 0;
	   enable = 0;
       baseAddr = 0;
       enableStore = 0;
       returnToBaseAddr = 0;
       incrementAddr = 0;
	end
	
	always begin
	   #2.5 clk = !clk;
	end

    always begin
        #5 samplePulse = !samplePulse;
    end
	
	task bitZero();
        begin
            dIn = 0;
            #10;
        end
    endtask
    task bitOne();
        begin
            dIn = 1;
            #10;
        end
    endtask

    task bigData();
        begin
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
        bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
        bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
            bitOne();
            bitOne();
            bitOne();
            bitZero();
            bitZero();
            bitOne();
        end
    endtask
    
    task increment();
        begin
            incrementAddr = 1;
            #20;
            incrementAddr = 0;
            #20;
        end
    endtask
    
    initial begin
        #25;
        resetN = 0;
        #45;
        resetN = 1;
        numFetches = 1;
        enableStore = 1;
        #5;
        enableStore = 0;
        #25
        enable = 1;
        #10;
        bigData();
        #40;
        enable = 0;
        #25;
        returnToBaseAddr = 1;
        #5;
        returnToBaseAddr = 0;
        #20;
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        #100;
        resetN = 0;
        #45;
        resetN = 1;
        baseAddr = 32'hC;
        numFetches = 1;
        enableStore = 1;
        #5;
        enableStore = 0;
        #25;
        returnToBaseAddr = 1;
        #5;
        returnToBaseAddr = 0;
        #20;
        enable = 1;
        #10;
        bigData();
        #40;
        enable = 0;
        #25;
        baseAddr = 0;
        numFetches = 1;
        enableStore = 1;
        #5;
        enableStore = 0;
        #25;
        returnToBaseAddr = 1;
        #5;
        returnToBaseAddr = 0;
        #20;
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        increment();
        #100;
    end
    

endmodule
